`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:32:14 11/08/2019 
// Design Name: 
// Module Name:    Semi_Procesador_64 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Semi_Procesador_64(
    input clk,
    input [7:0] SW,
    output [7:0] LEDS
    );
	 
	 


endmodule
